//------------------------------------------------------------------------------
//	Module:		Lab2Lock
//	Desc:			This module implements the functionality of a simple combination lock.
//					The lock uses 2 4-bit combination digits.
//					See the lab document for the suggested combination setting.
//	Params:		This module is not parameterized.
//	Inputs:		See Lab2 document
//	Outputs:	See Lab2 document
//
//	Author:     YOUR NAME GOES HERE
//------------------------------------------------------------------------------
module	Lab2Lock(
			//------------------------------------------------------------------
			//	Clock & Reset Inputs
			//------------------------------------------------------------------
			Clock,
			Reset,
			//------------------------------------------------------------------
			
			//------------------------------------------------------------------
			//	Inputs
			//------------------------------------------------------------------
			Enter,
			Digit,
			//------------------------------------------------------------------
			
			//------------------------------------------------------------------
			//	Outputs
			//------------------------------------------------------------------
			State,
			Open,
			Fail
			//------------------------------------------------------------------
	);
	//--------------------------------------------------------------------------
	//	Parameters
	//---------------------------------------
	localparam	DIGIT_1	=	4'h2,
					DIGIT_2	=	4'h3;
										
	//--------------------------------------------------------------------------
	
	//--------------------------------------------------------------------------
	//	Clock & Reset Inputs
	//--------------------------------------------------------------------------
	input					Clock;	// System clock
	input					Reset;	// System reset
	//--------------------------------------------------------------------------
	
	//--------------------------------------------------------------------------
	//	Inputs
	//--------------------------------------------------------------------------
	input					Enter;
	input		[3:0]		Digit;
	//--------------------------------------------------------------------------
	
	//--------------------------------------------------------------------------
	//	Outputs
	//--------------------------------------------------------------------------
	output		[2:0]		State;
	output		reg		Open;
	output		reg		Fail;
	//--------------------------------------------------------------------------

	//--------------------------------------------------------------------------
	//	State Encoding
	//--------------------------------------------------------------------------
	
	parameter LOCKED = 3'b000,
				 OK = 3'b001,
				 BAD1 = 3'b010,
				 BAD2 = 3'b011,
				 OPEN = 3'b100; 
	
	//--------------------------------------------------------------------------
	
	//--------------------------------------------------------------------------
	//	Wire Declarations
	//--------------------------------------------------------------------------
	
	reg [2:0] nome;
	
	//--------------------------------------------------------------------------
	
	//--------------------------------------------------------------------------
	//	Logic
	//--------------------------------------------------------------------------
	initial 
		nome = LOCKED;
	always @(posedge Clock && Reset) begin
		if (Reset)
			nome <= LOCKED;
		else begin
			case(nome) 
				LOCKED : begin
					if (Digit == DIGIT_1 && Enter)
						nome <= OK;
					else if(Enter)
						nome <= BAD1;
					Open = 0;
					Fail = 0;
				end
				OK : begin
					if (Digit == DIGIT_2 && Enter)
						nome <= OPEN;
					else if (Enter)
						nome <= BAD2;
					Open = 0;
					Fail = 0;
				end
				BAD1 : begin
					nome <= BAD2;
					Open = 0;
					Fail = 0;
				end
				BAD2 : begin
					nome <= BAD2;
					Open = 0;
					Fail = 1;
				end
				OPEN : begin
					Open = 1;
					Fail = 0;
				end
			endcase	
			end
	end
	
	assign State = nome;
	//--------------------------------------------------------------------------
endmodule
//------------------------------------------------------------------------------
